module tcgrom(addr, data);
  input [8:0] addr;
  output [7:0] data;
  reg [7:0] data;
  
  // A memory is implemented
  // using a case statement 
  
  always @(addr)
    begin
      case (addr)

        9'h008 : data = 8'b00011000; // %     **      %
        9'h009 : data = 8'b00111100; // %    ****     %
        9'h00a : data = 8'b01100110; // %   **  **    %
        9'h00b : data = 8'b01111110; // %   ******    %
        9'h00c : data = 8'b01100110; // %   **  **    %
        9'h00d : data = 8'b01100110; // %   **  **    %
        9'h00e : data = 8'b01100110; // %   **  **    %
        9'h00f : data = 8'b00000000; // %             %

        9'h018 : data = 8'b00111100; // %    ****     %
        9'h019 : data = 8'b01100110; // %   **  **    %
        9'h01a : data = 8'b01100000; // %   **        %
        9'h01b : data = 8'b01100000; // %   **        %
        9'h01c : data = 8'b01100000; // %   **        %
        9'h01d : data = 8'b01100110; // %   **  **    %
        9'h01e : data = 8'b00111100; // %    ****     %
        9'h01f : data = 8'b00000000; // %             %

        9'h028 : data = 8'b01111110; // %   ******    %
        9'h029 : data = 8'b01100000; // %   **        %
        9'h02a : data = 8'b01100000; // %   **        %
        9'h02b : data = 8'b01111000; // %   ****      %
        9'h02c : data = 8'b01100000; // %   **        %
        9'h02d : data = 8'b01100000; // %   **        %
        9'h02e : data = 8'b01111110; // %   ******    %
        9'h02f : data = 8'b00000000; // %             %


        9'h038 : data = 8'b00111100; // %    ****     %
        9'h039 : data = 8'b01100110; // %   **  **    %
        9'h03a : data = 8'b01100000; // %   **        %
        9'h03b : data = 8'b01101110; // %   ** ***    %
        9'h03c : data = 8'b01100110; // %   **  **    %
        9'h03d : data = 8'b01100110; // %   **  **    %
        9'h03e : data = 8'b00111100; // %    ****     %
        9'h03f : data = 8'b00000000; // %             %

        9'h040 : data = 8'b01100110; // %   **  **    %
        9'h041 : data = 8'b01100110; // %   **  **    %
        9'h042 : data = 8'b01100110; // %   **  **    %
        9'h043 : data = 8'b01111110; // %   ******    %
        9'h044 : data = 8'b01100110; // %   **  **    %
        9'h045 : data = 8'b01100110; // %   **  **    %
        9'h046 : data = 8'b01100110; // %   **  **    %
        9'h047 : data = 8'b00000000; // %             %

        9'h048 : data = 8'b00111100; // %    ****     %
        9'h049 : data = 8'b00011000; // %     **      %
        9'h04a : data = 8'b00011000; // %     **      %
        9'h04b : data = 8'b00011000; // %     **      %
        9'h04c : data = 8'b00011000; // %     **      %
        9'h04d : data = 8'b00011000; // %     **      %
        9'h04e : data = 8'b00111100; // %    ****     %
        9'h04f : data = 8'b00000000; // %             %

        9'h060 : data = 8'b01100000; // %   **        %
        9'h061 : data = 8'b01100000; // %   **        %
        9'h062 : data = 8'b01100000; // %   **        %
        9'h063 : data = 8'b01100000; // %   **        %
        9'h064 : data = 8'b01100000; // %   **        %
        9'h065 : data = 8'b01100000; // %   **        %
        9'h066 : data = 8'b01111110; // %   ******    %
        9'h067 : data = 8'b00000000; // %             %
	  
        9'h078 : data = 8'b00111100; // %    ****     %
        9'h079 : data = 8'b01100110; // %   **  **    %
        9'h07a : data = 8'b01100110; // %   **  **    %
        9'h07b : data = 8'b01100110; // %   **  **    %
        9'h07c : data = 8'b01100110; // %   **  **    %
        9'h07d : data = 8'b01100110; // %   **  **    %
        9'h07e : data = 8'b00111100; // %    ****     %
        9'h07f : data = 8'b00000000; // %             %

        9'h080 : data = 8'b01111100; // %   *****     %
        9'h081 : data = 8'b01100110; // %   **  **    %
        9'h082 : data = 8'b01100110; // %   **  **    %
        9'h083 : data = 8'b01111100; // %   *****     %
        9'h084 : data = 8'b01100000; // %   **        %
        9'h085 : data = 8'b01100000; // %   **        %
        9'h086 : data = 8'b01100000; // %   **        %
        9'h087 : data = 8'b00000000; // %             %

        9'h090 : data = 8'b01111100; // %   *****     %
        9'h091 : data = 8'b01100110; // %   **  **    %
        9'h092 : data = 8'b01100110; // %   **  **    %
        9'h093 : data = 8'b01111100; // %   *****     %
        9'h094 : data = 8'b01111000; // %   ****      %
        9'h095 : data = 8'b01101100; // %   ** **     %
        9'h096 : data = 8'b01100110; // %   **  **    %
        9'h097 : data = 8'b00000000; // %             %

        9'h098 : data = 8'b00111100; // %    ****     %
        9'h099 : data = 8'b01100110; // %   **  **    %
        9'h09a : data = 8'b01100000; // %   **        %
        9'h09b : data = 8'b00111100; // %    ****     %
        9'h09c : data = 8'b00000110; // %       **    %
        9'h09d : data = 8'b01100110; // %   **  **    %
        9'h09e : data = 8'b00111100; // %    ****     %
        9'h09f : data = 8'b00000000; // %             %

        9'h0a0 : data = 8'b01111110; // %   ******    %
        9'h0a1 : data = 8'b00011000; // %     **      %
        9'h0a2 : data = 8'b00011000; // %     **      %
        9'h0a3 : data = 8'b00011000; // %     **      %
        9'h0a4 : data = 8'b00011000; // %     **      %
        9'h0a5 : data = 8'b00011000; // %     **      %
        9'h0a6 : data = 8'b00011000; // %     **      %
        9'h0a7 : data = 8'b00000000; // %             %

        9'h0a8 : data = 8'b01100110; // %   **  **    %
        9'h0a9 : data = 8'b01100110; // %   **  **    %
        9'h0aa : data = 8'b01100110; // %   **  **    %
        9'h0ab : data = 8'b01100110; // %   **  **    %
        9'h0ac : data = 8'b01100110; // %   **  **    %
        9'h0ad : data = 8'b01100110; // %   **  **    %
        9'h0ae : data = 8'b00111100; // %    ****     %
        9'h0af : data = 8'b00000000; // %             %
 
 /*    
        9'h150 : data = 8'b00000000; // %             %
        9'h151 : data = 8'b01100110; // %   **  **    %
        9'h152 : data = 8'b00111100; // %    ****     %
        9'h153 : data = 8'b11111111; // %  ********   %
        9'h154 : data = 8'b00111100; // %    ****     %
        9'h155 : data = 8'b01100110; // %   **  **    %
        9'h156 : data = 8'b00000000; // %             %
        9'h157 : data = 8'b00000000; // %             %
*/

        9'h180 : data = 8'b00111100; // %    ****     %
        9'h181 : data = 8'b01100110; // %   **  **    %
        9'h182 : data = 8'b01101110; // %   ** ***    %
        9'h183 : data = 8'b01110110; // %   *** **    %
        9'h184 : data = 8'b01100110; // %   **  **    %
        9'h185 : data = 8'b01100110; // %   **  **    %
        9'h186 : data = 8'b00111100; // %    ****     %
        9'h187 : data = 8'b00000000; // %             %

        9'h188 : data = 8'b00011000; // %     **      %
        9'h189 : data = 8'b00011000; // %     **    . %
        9'h18a : data = 8'b00111000; // %    ***      %
        9'h18b : data = 8'b00011000; // %     **      %
        9'h18c : data = 8'b00011000; // %     **      %
        9'h18d : data = 8'b00011000; // %     **      %
        9'h18e : data = 8'b01111110; // %   ******    %
        9'h18f : data = 8'b00000000; // %             %

        9'h190 : data = 8'b00111100; // %    ****     %
        9'h191 : data = 8'b01100110; // %   **  **    %
        9'h192 : data = 8'b00000110; // %       **    %
        9'h193 : data = 8'b00001100; // %      **     %
        9'h194 : data = 8'b00110000; // %    **       %
        9'h195 : data = 8'b01100000; // %   **        %
        9'h196 : data = 8'b01111110; // %   ******    %
        9'h197 : data = 8'b00000000; // %             %

        9'h198 : data = 8'b00111100; // %    ****     %
        9'h199 : data = 8'b01100110; // %   **  **    %
        9'h19a : data = 8'b00000110; // %       **    %
        9'h19b : data = 8'b00011100; // %     ***     %
        9'h19c : data = 8'b00000110; // %       **    %
        9'h19d : data = 8'b01100110; // %   **  **    %
        9'h19e : data = 8'b00111100; // %    ****     %
        9'h19f : data = 8'b00000000; // %             %

        9'h1a0 : data = 8'b00000110; // %       **    %
        9'h1a1 : data = 8'b00001110; // %      ***    %
        9'h1a2 : data = 8'b00011110; // %     ****    %
        9'h1a3 : data = 8'b01100110; // %   **  **    %
        9'h1a4 : data = 8'b01111111; // %   *******   %
        9'h1a5 : data = 8'b00000110; // %       **    %
        9'h1a6 : data = 8'b00000110; // %       **    %
        9'h1a7 : data = 8'b00000000; // %             %

        9'h1a8 : data = 8'b01111110; // %   ******    %
        9'h1a9 : data = 8'b01100000; // %   **        %
        9'h1aa : data = 8'b01111100; // %   *****     %
        9'h1ab : data = 8'b00000110; // %       **    %
        9'h1ac : data = 8'b00000110; // %       **    %
        9'h1ad : data = 8'b01100110; // %   **  **    %
        9'h1ae : data = 8'b00111100; // %    ****     %
        9'h1af : data = 8'b00000000; // %             %

        9'h1b0 : data = 8'b00111100; // %    ****     %
        9'h1b1 : data = 8'b01100110; // %   **  **    %
        9'h1b2 : data = 8'b01100000; // %   **        %
        9'h1b3 : data = 8'b01111100; // %   *****     %
        9'h1b4 : data = 8'b01100110; // %   **  **    %
        9'h1b5 : data = 8'b01100110; // %   **  **    %
        9'h1b6 : data = 8'b00111100; // %    ****     %
        9'h1b7 : data = 8'b00000000; // %             %

        9'h1b8 : data = 8'b01111110; // %   ******    %
        9'h1b9 : data = 8'b01100110; // %   **  **    %
        9'h1ba : data = 8'b00001100; // %      **     %
        9'h1bb : data = 8'b00011000; // %     **      %
        9'h1bc : data = 8'b00011000; // %     **      %
        9'h1bd : data = 8'b00011000; // %     **      %
        9'h1be : data = 8'b00011000; // %     **      %
        9'h1bf : data = 8'b00000000; // %             %

        9'h1c0 : data = 8'b00111100; // %    ****     %
        9'h1c1 : data = 8'b01100110; // %   **  **    %
        9'h1c2 : data = 8'b01100110; // %   **  **    %
        9'h1c3 : data = 8'b00111100; // %    ****     %
        9'h1c4 : data = 8'b01100110; // %   **  **    %
        9'h1c5 : data = 8'b01100110; // %   **  **    %
        9'h1c6 : data = 8'b00111100; // %    ****     %
        9'h1c7 : data = 8'b00000000; // %             %

        9'h1c8 : data = 8'b00111100; // %    ****     %
        9'h1c9 : data = 8'b01100110; // %   **  **    %
        9'h1ca : data = 8'b01100110; // %   **  **    %
        9'h1cb : data = 8'b00111110; // %    *****    %
        9'h1cc : data = 8'b00000110; // %       **    %
        9'h1cd : data = 8'b01100110; // %   **  **    %
        9'h1ce : data = 8'b00111100; // %    ****     %
        9'h1cf : data = 8'b00000000; // %             %

	   //28
	   9'h0e0 : data = 8'b00011000; // %     **      %
        9'h0e1 : data = 8'b00011000; // %     **      %
        9'h0e2 : data = 8'b00011000; // %     **      %
        9'h0e3 : data = 8'b00011000; // %     **      %
        9'h0e4 : data = 8'b01111110; // %   ******    %
        9'h0e5 : data = 8'b00111100; // %    ****     %
        9'h0e6 : data = 8'b00011000; // %     **      %
        9'h0e7 : data = 8'b00000000; // %             %

	   //29
        9'h0e8 : data = 8'b00000000; // %    ****     %
        9'h0e9 : data = 8'b00010000; // %      **     %
        9'h0ea : data = 8'b00011000; // %      **     %
        9'h0eb : data = 8'b01111110; // %      **     %
        9'h0ec : data = 8'b01111110; // %      **     %
        9'h0ed : data = 8'b00011000; // %      **     %
        9'h0ee : data = 8'b00010000; // %    ****     %
        9'h0ef : data = 8'b00000000; // %             %

	   //30
        9'h0f0 : data = 8'b00000000; // %             %
        9'h0f1 : data = 8'b00011000; // %     **      %
        9'h0f2 : data = 8'b00111100; // %    ****     %
        9'h0f3 : data = 8'b01111110; // %   ******    %
        9'h0f4 : data = 8'b00011000; // %     **      %
        9'h0f5 : data = 8'b00011000; // %     **      %
        9'h0f6 : data = 8'b00011000; // %     **      %
        9'h0f7 : data = 8'b00011000; // %     **      %

	   //31
        9'h0f8 : data = 8'b00000000; // %             %
        9'h0f9 : data = 8'b00010000; // %     *       %
        9'h0fa : data = 8'b00110000; // %    **       %
        9'h0fb : data = 8'b01111111; // %   *******   %
        9'h0fc : data = 8'b01111111; // %   *******   %
        9'h0fd : data = 8'b00110000; // %    **       %
        9'h0fe : data = 8'b00010000; // %     *       %
        9'h0ff : data = 8'b00000000; // %             %


		default: data = 8'd0;
      endcase
    end

endmodule
