module score();



endmodule
